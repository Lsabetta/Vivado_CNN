library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
use work.fixed_generic_pkg.all;
use work.fixed_float_types.all;
use work.my_types.all;

package my_weights is

  constant w_1: matrix9 := ((to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits)),
                            (to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits)),
                            (to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits)));

  constant b_1: thresholds_conv1 := (others => to_sfixed(0.375, w_ibits, w_fbits));

  constant w_2: matrix9 := ((to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits)),
                            (to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits)),
                            (to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits)));

  constant b_2: thresholds_conv1 := (others => to_sfixed(0.25, w_ibits, w_fbits));

  constant w_3: matrix6_9 := (((to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits)),
                              (to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits)),
                              (to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits))),

                              ((to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits)),
                              (to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits)),
                              (to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits))),

                              ((to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits)),
                              (to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits)),
                              (to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits))),

                              ((to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits)),
                              (to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits)),
                              (to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits))),

                              ((to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits)),
                              (to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits)),
                              (to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits))),

                              ((to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits)),
                              (to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits)),
                              (to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits))));

  constant b_3: thresholds_conv6 := (to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits));

  constant w_4: matrix6_9_6 := ((((to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits)),
                                (to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits)),
                                (to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits))),
                                ((to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits)),
                                (to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits)),
                                (to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits))),
                                ((to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits)),
                                (to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits)),
                                (to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits)))),

                                (((to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits)),
                                (to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits)),
                                (to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits))),
                                ((to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits)),
                                (to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits)),
                                (to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits))),
                                ((to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits)),
                                (to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits)),
                                (to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits)))),

                                (((to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits)),
                                (to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits)),
                                (to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits))),
                                ((to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits)),
                                (to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits)),
                                (to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits))),
                                ((to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits)),
                                (to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits)),
                                (to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits)))),

                                (((to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits)),
                                (to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits)),
                                (to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits))),
                                ((to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits)),
                                (to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits)),
                                (to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits))),
                                ((to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits)),
                                (to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits)),
                                (to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits)))),

                                (((to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits)),
                                (to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits)),
                                (to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits))),
                                ((to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits)),
                                (to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits)),
                                (to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits))),
                                ((to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits)),
                                (to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits)),
                                (to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits)))),

                                (((to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits)),
                                (to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits)),
                                (to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits))),
                                ((to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits)),
                                (to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits)),
                                (to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits))),
                                ((to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits)),
                                (to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits)),
                                (to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits)))));

  constant b_4: thresholds_conv6 := (to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits));

  constant dw_1: matrix10_48 := ((to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits)),
                                 (to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits)),
                                 (to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits)),
                                 (to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits)),
                                 (to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits)),
                                 (to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits)),
                                 (to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits)),
                                 (to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits)),
                                 (to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits)),
                                 (to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits)));

  constant db_1: thresholds_dense := (to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits));

  constant dw_2: matrix10_10 := ((to_sfixed(-0.3125, w_ibits, w_fbits), to_sfixed(-0.1875, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.0625, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.4375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.0625, w_ibits, w_fbits), to_sfixed(-0.3125, w_ibits, w_fbits)),
                                 (to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits)),
                                 (to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits)),
                                 (to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits)),
                                 (to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits)),
                                 (to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.75, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.625, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.75, w_ibits, w_fbits)),
                                 (to_sfixed(0.75, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.5, w_ibits, w_fbits), to_sfixed(0.875, w_ibits, w_fbits)),
                                 (to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(0.25, w_ibits, w_fbits), to_sfixed(-0.625, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits)),
                                 (to_sfixed(-0.1875, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.1875, w_ibits, w_fbits), to_sfixed(-0.1875, w_ibits, w_fbits), to_sfixed(0.4375, w_ibits, w_fbits), to_sfixed(0.375, w_ibits, w_fbits), to_sfixed(0.0625, w_ibits, w_fbits), to_sfixed(-0.1875, w_ibits, w_fbits), to_sfixed(0.4375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits)),
                                 (to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.0, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(-0.875, w_ibits, w_fbits), to_sfixed(-0.5, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits)));

  constant db_2: thresholds_dense := (to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(-0.125, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.375, w_ibits, w_fbits), to_sfixed(0.125, w_ibits, w_fbits), to_sfixed(-0.25, w_ibits, w_fbits));

  constant dw_3: matrix2_10 := ((to_sfixed(0.021518826, w_ibits_out, w_fbits_out), to_sfixed(0.069911405, w_ibits_out, w_fbits_out), to_sfixed(-0.1881477, w_ibits_out, w_fbits_out), to_sfixed(0.1553226, w_ibits_out, w_fbits_out), to_sfixed(-0.0042044595, w_ibits_out, w_fbits_out), to_sfixed(0.24569526, w_ibits_out, w_fbits_out), to_sfixed(0.26121324, w_ibits_out, w_fbits_out), to_sfixed(-0.22705604, w_ibits_out, w_fbits_out), to_sfixed(-0.057761535, w_ibits_out, w_fbits_out), to_sfixed(-0.27830175, w_ibits_out, w_fbits_out)),
                                (to_sfixed(-0.6931504, w_ibits_out, w_fbits_out), to_sfixed(0.007868746, w_ibits_out, w_fbits_out), to_sfixed(-0.0400587, w_ibits_out, w_fbits_out), to_sfixed(0.009778387, w_ibits_out, w_fbits_out), to_sfixed(-0.041952062, w_ibits_out, w_fbits_out), to_sfixed(0.00067524565, w_ibits_out, w_fbits_out), to_sfixed(0.0072312234, w_ibits_out, w_fbits_out), to_sfixed(-0.015551189, w_ibits_out, w_fbits_out), to_sfixed(0.011560225, w_ibits_out, w_fbits_out), to_sfixed(-0.03564694, w_ibits_out, w_fbits_out)));

  constant db_3: thresholds_out := (to_sfixed(0.22447677, w_ibits_out, w_fbits_out), to_sfixed(0.50014687, w_ibits_out, w_fbits_out));














end package;
